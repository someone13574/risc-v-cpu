module control_unit(
    input clk,
    input logic clk_enable,
    input [31:0] microcode_s0,
    input [24:0] instruction_data_s0,
    input [29:0] jump_location,
    input [31:0] reg_out_a,
    input [31:0] reg_out_b,
    output reg [29:0] pc,
    output reg [29:0] pc_s2,
    output reg [24:0] instruction_data_s3,
    output [3:0] alu_op_select,
    output pre_alu_a_to_alu_a,
    output [1:0] pre_alu_a_select,
    output pre_alu_b_to_alu_b,
    output [1:0] pre_alu_b_select,
    output mem_we,
    output alu_out_to_mem_addr,
    output reg_we,
    output up_to_reg_data_in,
    output alu_out_to_reg_data_in,
    output ret_addr_to_reg_data_in,
    output mem_data_to_reg_data_in,
    output block_inst,
    output reg [31:0] microcode_s1,
    output reg [31:0] microcode_s2,
    output reg [31:0] microcode_s3
);

typedef enum bit[2:0] {
    NULL_CMP_OP        = 3'b000,
    EQ_CMP_OP          = 3'b001,
    NOT_EQ_CMP_OP      = 3'b010,
    LESS_THAN_CMP_OP   = 3'b011,
    GREATER_EQ_CMP_OP  = 3'b100,
    LESS_THAN_U_CMP_OP = 3'b101,
    GREATER_EQ_U_CM_OP = 3'b110,
    TRUE_CMP_OP        = 3'b111
} cmp_ops_e;

reg [29:0] pc_si;
reg [29:0] pc_s0;
reg [29:0] pc_s1;

// reg [31:0] microcode_s1;
// reg [31:0] microcode_s2;
// reg [31:0] microcode_s3;

reg [24:0] instruction_data_s1;
reg [24:0] instruction_data_s2;

reg branch;
wire jump_if_branch;
wire data_dep_with_s1;
wire data_dep_with_s2;
wire data_dep_with_s3;
wire data_dep;

reg hold;
reg [24:0] held_instruction_data;

assign data_dep_with_s1 = (((rs1_s0 == rd_s1) & check_rs1_dep) | ((rs2_s0 == rd_s1) & check_rs2_dep)) & reg_we_s1;
assign data_dep_with_s2 = (((rs1_s0 == rd_s2) & check_rs1_dep) | ((rs2_s0 == rd_s2) & check_rs2_dep)) & reg_we_s2;
assign data_dep_with_s3 = (((rs1_s0 == rd_s3) & check_rs1_dep) | ((rs2_s0 == rd_s3) & check_rs2_dep)) & reg_we;
assign data_dep = data_dep_with_s1 | data_dep_with_s2 | data_dep_with_s3;

wire block_for_branch = microcode_s0[17] | microcode_s1[17] | microcode_s2[17] | microcode_s3[17]; // jump if branch mc
wire mem_in_use;
wire mem_in_use_s3;
assign block_inst = mem_in_use_s3 | data_dep | hold | block_for_branch;

wire [2:0] branch_cond_select;
always @(posedge clk) begin
    if (clk_enable) begin
        if (jump_if_branch & branch) begin
            pc <= jump_location;
        end else if (data_dep) begin
            pc <= pc_s0;
        end else if (hold & mem_in_use) begin
            pc <= pc_s1;
        end else if (mem_in_use) begin
            pc <= pc_si;
        end else begin
            pc <= pc + 30'b1;
        end

        hold <= data_dep;

        case (branch_cond_select)
            NULL_CMP_OP:        branch <= 1'b0;
            EQ_CMP_OP:          branch <= reg_out_a          == reg_out_b;
            NOT_EQ_CMP_OP:      branch <= reg_out_a          != reg_out_b;
            LESS_THAN_CMP_OP:   branch <= $signed(reg_out_a) <  $signed(reg_out_b);
            GREATER_EQ_CMP_OP:  branch <= $signed(reg_out_a) >= $signed(reg_out_b);
            LESS_THAN_U_CMP_OP: branch <= reg_out_a          <  reg_out_b;
            GREATER_EQ_U_CM_OP: branch <= reg_out_a          >= reg_out_b;
            TRUE_CMP_OP:        branch <= 1'b1;
        endcase

        pc_si <= pc;
        pc_s0 <= pc_si;
        pc_s1 <= pc_s0;
        pc_s2 <= pc_s1;

        microcode_s1 <= (data_dep) ? 32'b00000000 : microcode_s0;
        microcode_s2 <= microcode_s1;
        microcode_s3 <= microcode_s2;

        instruction_data_s1 <= instruction_data_s0;
        instruction_data_s2 <= instruction_data_s1;
        instruction_data_s3 <= instruction_data_s2;
    end
end

// s0 signals
wire check_rs1_dep = microcode_s0[0];
wire check_rs2_dep = microcode_s0[1];
assign pre_alu_a_select = microcode_s0[3:2];
assign pre_alu_b_select = microcode_s0[5:4];

// s1 signals
assign pre_alu_a_to_alu_a = microcode_s1[6];
assign pre_alu_b_to_alu_b = microcode_s1[7];
assign alu_op_select      = microcode_s1[11:8];
assign branch_cond_select = microcode_s1[14:12];

// s2 signals
assign mem_we                = microcode_s2[15];
assign alu_out_to_mem_addr   = microcode_s2[16];
assign jump_if_branch        = microcode_s2[17];
assign mem_in_use            = microcode_s2[18];

// s3 signals
assign mem_in_use_s3           = microcode_s3[18];
assign reg_we                  = microcode_s3[19]; // update reg_we_s1 & reg_we_s2 as well
assign up_to_reg_data_in       = microcode_s3[20];
assign alu_out_to_reg_data_in  = microcode_s3[21];
assign ret_addr_to_reg_data_in = microcode_s3[22];
assign mem_data_to_reg_data_in = microcode_s3[23];

// data dep signals (s1, s2)
wire reg_we_s1 = microcode_s1[19];
wire reg_we_s2 = microcode_s2[19];

wire [4:0] rs1_s0 = instruction_data_s0[12:8];
wire [4:0] rs2_s0 = instruction_data_s0[17:13];

wire [4:0] rd_s1 = instruction_data_s1[4:0];
wire [4:0] rd_s2 = instruction_data_s2[4:0];
wire [4:0] rd_s3 = instruction_data_s3[4:0];

endmodule

// si = first stage with decoded instruction
// s0 = read
// s1 = execute
// s2 = read/write memory & pc
// s3 = write regs
