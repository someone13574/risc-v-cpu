module risc_v_core(
	input clk
);



endmodule